package pack1;
import uvm_pkg::*;
`include "uvm_macros.svh"
`include "seq_item.svh"
`include "sequence.svh"
`include "driver.svh"
`include "monitor.svh"
`include "sequencer.svh"
`include "agent.svh"
`include "scoreboard.svh"
`include "subscriber.svh"
`include "env.svh"
`include "test.svh"
endpackage