package pack;
  `include "Trans.svh"
  `include "Sequencer.svh"
  `include "Driver.svh"
  `include "Monitor.svh"
  `include "Scoreboard.svh"
  `include "Subscriber.svh"
  `include "Env.svh"
endpackage
